* SPICE netlist written by S-Edit Win32 6.00
* Written on Jan 14, 2024 at 01:05:09

* Waveform probing commands
.probe
.options probefilename="FA1bit"
+ probesdbfile="X:\Q2_S_edit\FA1bit.sdb"
+ probetopmodule="Addr_8bit"

* No Ports in cell: PageID_Tanner
* End of module with no ports: PageID_Tanner

.SUBCKT XOR2 A B Out Gnd Vdd
M1 N2 B Gnd Gnd NMOS W='22*l' L='2*l' AS='66*l*l' AD='66*l*l' PS='24*l' PD='24*l' M=1
M2 N2 A Gnd Gnd NMOS W='22*l' L='2*l' AS='66*l*l' AD='66*l*l' PS='24*l' PD='24*l' M=1
M6 Out B N3 Gnd NMOS W='22*l' L='2*l' AS='66*l*l' AD='66*l*l' PS='24*l' PD='24*l' M=1
M5 N3 A Gnd Gnd NMOS W='22*l' L='2*l' AS='66*l*l' AD='66*l*l' PS='24*l' PD='24*l' M=1
M9 Out N2 Gnd Gnd NMOS W='22*l' L='2*l' AS='66*l*l' AD='66*l*l' PS='24*l' PD='24*l' M=1
* Page Size:  5x7
* S-Edit  2-Input XOR Gate (TIB)
* Designed by: J. Luo  Jan 14, 2024  00:50:24
* Schematic generated by S-Edit
* from file X:\Q2_S_edit\FA1bit / module XOR2 / page Page0 
M3 N2 B N6 Vdd PMOS W='22*l' L='2*l' AS='66*l*l' AD='66*l*l' PS='24*l' PD='24*l' M=1
M4 N6 A Vdd Vdd PMOS W='22*l' L='2*l' AS='66*l*l' AD='66*l*l' PS='24*l' PD='24*l' M=1
M7 N5 A Vdd Vdd PMOS W='22*l' L='2*l' AS='66*l*l' AD='66*l*l' PS='24*l' PD='24*l' M=1
M10B Out N2 N5 Vdd PMOS W='22*l' L='2*l' AS='66*l*l' AD='66*l*l' PS='24*l' PD='24*l' M=1
M8 N4 B Vdd Vdd PMOS W='22*l' L='2*l' AS='66*l*l' AD='66*l*l' PS='24*l' PD='24*l' M=1
M10 Out N2 N4 Vdd PMOS W='22*l' L='2*l' AS='66*l*l' AD='66*l*l' PS='24*l' PD='24*l' M=1
.ENDS

.SUBCKT NAND2 A B Out Gnd Vdd
M3 Out B 1 Gnd NMOS W='28*l' L='2*l' AS='148*l*l' AD='84*l*l' PS='68*l' PD='34*l' M=1
M4 1 A Gnd Gnd NMOS W='28*l' L='2*l' AS='84*l*l' AD='144*l*l' PS='34*l' PD='68*l' M=1
* Page Size:  5x7
* S-Edit  2-Input NAND Gate (TIB)
* Designed by: J. Luo  Jan 14, 2024  00:50:24
* Schematic generated by S-Edit
* from file X:\Q2_S_edit\FA1bit / module NAND2 / page Page0 
M2 Out B Vdd Vdd PMOS W='28*l' L='2*l' AS='144*l*l' AD='84*l*l' PS='68*l' PD='34*l' M=1
M1 Out A Vdd Vdd PMOS W='28*l' L='2*l' AS='84*l*l' AD='144*l*l' PS='34*l' PD='68*l' M=1
.ENDS

.SUBCKT FA1bit A B Cin Cout Sum Gnd Vdd
XNAND2_3 Cin N9 N6 Gnd Vdd NAND2
XNAND2_4 N6 N13 Cout Gnd Vdd NAND2
XNAND2_5 B A N13 Gnd Vdd NAND2
XXOR2_1 A B N9 Gnd Vdd XOR2
XXOR2_2 N9 Cin Sum Gnd Vdd XOR2
.ENDS

.SUBCKT Pad_Bond SIGNAL Subs
C1 SIGNAL Subs 0.25pF
* Page Size:  5x7
* S-Edit  Output Pad
* Designed by: D.Gunawan, J.Luo, K.Schaefer  Jan 14, 2024  00:55:10
* Schematic generated by S-Edit
* from file X:\Q2_S_edit\FA1bit / module Pad_Bond / page Page0 
.ENDS

.SUBCKT PadBidirHE_2.0u DataIn DataInB DataInUnBuf DataOut OE Pad Gnd Subs Vdd
MN_4_1 OEB OE Gnd Gnd NMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=1
MN_4_2 N29 DataOut Gnd Gnd NMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=1
MN_4_3 N20 OE N29 Gnd NMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=1
MN_4_4 N29 OEB Gnd Gnd NMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=1
MN_4_5 Pad N29 Gnd Gnd NMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=10
MN_4_6 DataInB DataInUnBuf Gnd Gnd NMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=2
MN_4_7 DataIn DataInB Gnd Gnd NMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=4
XPad_Bond_1 Pad Subs Pad_Bond
* Page Size:  5x7
* S-Edit  Bidirectional Pad
* Designed by: D.Gunawan, J.Luo  Jan 14, 2024  00:55:10
* Schematic generated by S-Edit
* from file X:\Q2_S_edit\FA1bit / module PadBidirHE_2.0u / page Page0 
MP_4_1 OEB OE Vdd Vdd PMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=1
MP_4_2 N20 DataOut Vdd Vdd PMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=2
MP_4_3 N29 OEB N20 Vdd PMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=2
MP_4_4 N20 OE Vdd Vdd PMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=1
MP_4_5 Pad N20 Vdd Vdd PMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=10
MP_4_6 DataInB DataInUnBuf Vdd Vdd PMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=2
MP_4_7 DataIn DataInB Vdd Vdd PMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=4
R1 Pad DataInUnBuf 100 TC1=0.0 TC2=0.0
.ENDS

.SUBCKT PadBidirHE DataIn DataInB DataInUnBuf DataOut OE Pad Gnd Subs Vdd
XPadBidirHE_2.0u_1 DataIn DataInB DataInUnBuf DataOut OE Pad Gnd Subs Vdd
+ PadBidirHE_2.0u
* Page Size:  5x7
* S-Edit  Bidirectional Pad
* Designed by: D.Gunawan, J.Luo  Jan 14, 2024  00:55:10
* Schematic generated by S-Edit
* from file X:\Q2_S_edit\FA1bit / module PadBidirHE / page Page0 
.ENDS

.SUBCKT PadInC DataIn DataInB DataInUnBuf Pad Gnd Subs Vdd
XPadBidirHE_1 DataIn DataInB DataInUnBuf Gnd Gnd Pad Gnd Subs Vdd PadBidirHE
* Page Size:  5x7
* S-Edit  Input Pad
* Designed by: D.Gunawan, J.Luo  Jan 14, 2024  00:52:34
* Schematic generated by S-Edit
* from file X:\Q2_S_edit\FA1bit / module PadInC / page Page0 
.ENDS

.SUBCKT PadOut DataOut Pad Gnd Subs Vdd
XPadBidirHE_1 N6 N5 N4 DataOut Vdd Pad Gnd Subs Vdd PadBidirHE
* Page Size:  5x7
* S-Edit  Output Pad
* Designed by: D.Gunawan, J.Luo  Jan 14, 2024  00:55:10
* Schematic generated by S-Edit
* from file X:\Q2_S_edit\FA1bit / module PadOut / page Page0 
.ENDS

* Main circuit: Addr_8bit
XFA1bit_1 N1 N2 N3 N8 N5 Gnd Vdd FA1bit
XFA1bit_2 N6 N7 N8 N13 N10 Gnd Vdd FA1bit
XFA1bit_3 N11 N12 N13 N18 N15 Gnd Vdd FA1bit
XFA1bit_4 N16 N17 N18 N23 N20 Gnd Vdd FA1bit
XFA1bit_5 N21 N22 N23 N28 N25 Gnd Vdd FA1bit
XFA1bit_6 N26 N27 N28 N33 N30 Gnd Vdd FA1bit
XFA1bit_7 N31 N32 N33 N38 N35 Gnd Vdd FA1bit
XFA1bit_8 N36 N37 N38 N39 N40 Gnd Vdd FA1bit
XPadInC_1 N1 N43 N42 a0 Gnd Subs Vdd PadInC
XPadInC_2 N2 N46 N45 b0 Gnd Subs Vdd PadInC
XPadInC_3 N6 N49 N48 a1 Gnd Subs Vdd PadInC
XPadInC_4 N7 N52 N51 b1 Gnd Subs Vdd PadInC
XPadInC_5 N11 N55 N54 a2 Gnd Subs Vdd PadInC
XPadInC_6 N12 N58 N57 b2 Gnd Subs Vdd PadInC
XPadInC_7 N16 N61 N60 a3 Gnd Subs Vdd PadInC
XPadInC_8 N17 N64 N63 b3 Gnd Subs Vdd PadInC
XPadInC_9 N21 N67 N66 a4 Gnd Subs Vdd PadInC
XPadInC_10 N22 N70 N69 b4 Gnd Subs Vdd PadInC
XPadInC_11 N26 N73 N72 a5 Gnd Subs Vdd PadInC
XPadInC_12 N27 N76 N75 b5 Gnd Subs Vdd PadInC
XPadInC_13 N31 N79 N78 a6 Gnd Subs Vdd PadInC
XPadInC_14 N32 N82 N81 b6 Gnd Subs Vdd PadInC
XPadInC_15 N36 N85 N84 a7 Gnd Subs Vdd PadInC
XPadInC_16 N37 N88 N87 b7 Gnd Subs Vdd PadInC
XPadInC_17 N3 N91 N90 Cin Gnd Subs Vdd PadInC
XPadOut_1 N5 Sum0 Gnd Subs Vdd PadOut
XPadOut_2 N10 Sum1 Gnd Subs Vdd PadOut
XPadOut_3 N15 Sum2 Gnd Subs Vdd PadOut
XPadOut_4 N20 Sum3 Gnd Subs Vdd PadOut
XPadOut_5 N25 Sum4 Gnd Subs Vdd PadOut
XPadOut_6 N30 Sum5 Gnd Subs Vdd PadOut
XPadOut_7 N35 Sum6 Gnd Subs Vdd PadOut
XPadOut_8 N40 Sum7 Gnd Subs Vdd PadOut
XPadOut_9 N39 Cout Gnd Subs Vdd PadOut
* End of main circuit: Addr_8bit
